package testbench_pkg;

parameter CLOCK_SPEED = 50; // 10MHZ
parameter TB_TIME_OUT_MS = 1; // testbench timeout in miliseconds

endpackage