../../../utils/utils.sv