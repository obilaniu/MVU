/**
 * Vector-Vector Product.
 */


/**** Module vvp ****/
module vvp(mode, W, D, S);


/* Parameters */
parameter  n  = 64;

localparam a  = $clog2(n);
localparam nr = (1 << a)/2;
localparam nl = n-nr;
localparam ar = $clog2(nr);
localparam al = $clog2(nl);

input  wire[     1 : 0] mode;
input  wire[   n-1 : 0] W;
input  wire[ 2*n-1 : 0] D;

output wire[ a+2-1 : 0] S;


/* Locals */
wire       [ar+2-1 : 0] Sr;
wire       [al+2-1 : 0] Sl;


/* Modal Multiplier Logic */
function [1:0] vvp_func(input[1:0] fmode,
                        input[0:0] fW,
                        input[1:0] fD);
begin
	if         (fmode == 2'b00) begin /* Weights {+1,-1} */
		vvp_func = fW ?   -fD :   +fD;
	end else if(fmode == 2'b01) begin /* Weights { 0,+1} */
		vvp_func = fW ?   +fD : 2'b00;
	end else if(fmode == 2'b10) begin /* Weights { 0,-1} */
		vvp_func = fW ?   -fD : 2'b00;
	end else                    begin /* Weights { 0, 0} */
		vvp_func = fW ? 2'b00 : 2'b00;
	end
end
endfunction


/* Recursive Hardware Logic Generation */
generate if(n == 1) begin
	assign S = vvp_func(mode, W, D);
end else if(n >= 2) begin
	vvp #(nr) r (mode, W[ 0 +: nr], D[  0  +: 2*nr], Sr);
	vvp #(nl) l (mode, W[nr +: nl], D[2*nr +: 2*nl], Sl);
	assign S = {{(a-al){Sl[al+1]}}, Sl} + {{(a-ar){Sr[ar+1]}}, Sr};
end endgenerate


/* Module end */
endmodule





/**** Test Module test_vvp ****/
module test_vvp();


/* Local parameters for test */
localparam n = 64;
localparam a = $clog2(n);


/* Create input registers and output wires */
reg        [    1 : 0] mode;
reg        [  n-1 : 0] W;
reg  signed[2*n-1 : 0] D;
wire signed[a+2-1 : 0] S;


/* Create instance */
vvp #(n) master (mode, W, D, S);


/* Run test */
initial begin
	$display("Testing %1d-wide Vector-Vector Dot Product...", n);
	$display("Testing Mode 00 {+1,-1} ...");
	assign mode = 2'b00;
	assign W = {n{ 1'b0}};
	assign D = {n{-2'd1}}; #1; $display("+1 * -1 = -1 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display("+1 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display("+1 * +1 =  1 ? %d", S); #1;
	assign W = {n{ 1'b1}};
	assign D = {n{-2'd1}}; #1; $display("-1 * -1 =  1 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display("-1 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display("-1 * +1 = -1 ? %d", S); #1;
	
	$display("Testing Mode 01 { 0,+1} ...");
	assign mode = 2'b01;
	assign W = {n{ 1'b0}};
	assign D = {n{-2'd1}}; #1; $display(" 0 * -1 =  0 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display(" 0 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display(" 0 * +1 =  0 ? %d", S); #1;
	assign W = {n{ 1'b1}};
	assign D = {n{-2'd1}}; #1; $display("+1 * -1 = -1 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display("+1 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display("+1 * +1 =  1 ? %d", S); #1;
	
	$display("Testing Mode 10 { 0,-1} ...");
	assign mode = 2'b10;
	assign W = {n{ 1'b0}};
	assign D = {n{-2'd1}}; #1; $display(" 0 * -1 =  0 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display(" 0 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display(" 0 * +1 =  0 ? %d", S); #1;
	assign W = {n{ 1'b1}};
	assign D = {n{-2'd1}}; #1; $display("-1 * -1 =  1 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display("-1 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display("-1 * +1 = -1 ? %d", S); #1;
	
	$display("Testing Mode 11 { 0, 0} ...");
	assign mode = 2'b11;
	assign W = {n{ 1'b0}};
	assign D = {n{-2'd1}}; #1; $display(" 0 * -1 =  0 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display(" 0 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display(" 0 * +1 =  0 ? %d", S); #1;
	assign W = {n{ 1'b1}};
	assign D = {n{-2'd1}}; #1; $display(" 0 * -1 =  0 ? %d", S); #1;
	assign D = {n{+2'd0}}; #1; $display(" 0 *  0 =  0 ? %d", S); #1;
	assign D = {n{+2'd1}}; #1; $display(" 0 * +1 =  0 ? %d", S); #1;
	
	$display("");
	assign mode = 2'b00;
	assign W = {n{ 1'b0}};
	assign D = {n{-2'b1}};
	#1;
	$display("mode = '%b'", mode);
	$display("W    = '%b'", W);
	$display("D    = '%b'", D);
	$display("master.Sr = '%b'", master.Sr);
	$display("master.Sl = '%b'", master.Sl);
	$display("master.S  = '%b'", master.S);
	$display("S    = '%d'", S);
end

endmodule
