//================================================================
// Simulation macros
//================================================================

//================================================================
// hard coded HDL paths for verification 
//================================================================
