module toplevel();

initial begin
	
end

endmodule
